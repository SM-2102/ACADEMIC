module notgate(input a, output b);
  assign b = ~a;
endmodule
